`include "APB_DEFINE.sv"
`include "APB_INTERFACE.sv"
package pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;
`include "APB_TRANS.sv"
`include "APB_SEQUENCE.sv"
`include "APB_SEQUENCER.sv"
`include "APB_DRIVER.sv"
`include "APB_MONITOR.sv"
`include "APB_AGENT.sv"
`include "APB_reference_model.sv"
`include "APB_SCOREBOARD.sv"
`include "APB_ENV.sv"
`include "APB_TEST.sv"

endpackage
